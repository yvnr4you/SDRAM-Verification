/////////////////////////////////////////////////////////////////
////        This is the package file.                        ////
////                                                         ////
////                                                         ////
////     Created By: Manasa Gurrala                          ////
////                 Venkata Naveen Reddy Yalla              ////
////                 Karthik Rudraraju                       ////
////                                                         ////
/////////////////////////////////////////////////////////////////

package sdrctrl_package;
import uvm_pkg::*;

`include "uvm_macros.svh"
`include "coverage.svh"
`include "stimulus_tester.svh"
`include "stimulus_values.svh"
`include "scoreboard.svh"
`include "env.svh"
`include "test.svh"


endpackage : sdrctrl_package
